sync_sync_out_altiobuf_inst : sync_sync_out_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
