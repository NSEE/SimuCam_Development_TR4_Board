spwc_spw_rx_altiobuf_inst : spwc_spw_rx_altiobuf PORT MAP (
		datain	 => datain_sig,
		datain_b	 => datain_b_sig,
		dataout	 => dataout_sig
	);
