-- MebX_Qsys_Project.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project is
	port (
		board_led_export                                            : out   std_logic_vector(3 downto 0);                     --                            board_led.export
		button_export                                               : in    std_logic_vector(3 downto 0)  := (others => '0'); --                               button.export
		clk50_clk                                                   : in    std_logic                     := '0';             --                                clk50.clk
		csense_adc_fo_export                                        : out   std_logic;                                        --                        csense_adc_fo.export
		csense_cs_n_export                                          : out   std_logic_vector(1 downto 0);                     --                          csense_cs_n.export
		csense_sck_export                                           : out   std_logic;                                        --                           csense_sck.export
		csense_sdi_export                                           : out   std_logic;                                        --                           csense_sdi.export
		csense_sdo_export                                           : in    std_logic                     := '0';             --                           csense_sdo.export
		m0_ddr3_i2c_scl_export                                      : out   std_logic;                                        --                      m0_ddr3_i2c_scl.export
		m0_ddr3_i2c_sda_export                                      : inout std_logic                     := '0';             --                      m0_ddr3_i2c_sda.export
		m0_ddr3_memory_mem_a                                        : out   std_logic_vector(13 downto 0);                    --                       m0_ddr3_memory.mem_a
		m0_ddr3_memory_mem_ba                                       : out   std_logic_vector(2 downto 0);                     --                                     .mem_ba
		m0_ddr3_memory_mem_ck                                       : out   std_logic_vector(0 downto 0);                     --                                     .mem_ck
		m0_ddr3_memory_mem_ck_n                                     : out   std_logic_vector(0 downto 0);                     --                                     .mem_ck_n
		m0_ddr3_memory_mem_cke                                      : out   std_logic_vector(0 downto 0);                     --                                     .mem_cke
		m0_ddr3_memory_mem_cs_n                                     : out   std_logic_vector(0 downto 0);                     --                                     .mem_cs_n
		m0_ddr3_memory_mem_dm                                       : out   std_logic_vector(7 downto 0);                     --                                     .mem_dm
		m0_ddr3_memory_mem_ras_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_ras_n
		m0_ddr3_memory_mem_cas_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_cas_n
		m0_ddr3_memory_mem_we_n                                     : out   std_logic_vector(0 downto 0);                     --                                     .mem_we_n
		m0_ddr3_memory_mem_reset_n                                  : out   std_logic;                                        --                                     .mem_reset_n
		m0_ddr3_memory_mem_dq                                       : inout std_logic_vector(63 downto 0) := (others => '0'); --                                     .mem_dq
		m0_ddr3_memory_mem_dqs                                      : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs
		m0_ddr3_memory_mem_dqs_n                                    : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs_n
		m0_ddr3_memory_mem_odt                                      : out   std_logic_vector(0 downto 0);                     --                                     .mem_odt
		m0_ddr3_memory_pll_sharing_pll_mem_clk                      : out   std_logic;                                        --           m0_ddr3_memory_pll_sharing.pll_mem_clk
		m0_ddr3_memory_pll_sharing_pll_write_clk                    : out   std_logic;                                        --                                     .pll_write_clk
		m0_ddr3_memory_pll_sharing_pll_locked                       : out   std_logic;                                        --                                     .pll_locked
		m0_ddr3_memory_pll_sharing_pll_write_clk_pre_phy_clk        : out   std_logic;                                        --                                     .pll_write_clk_pre_phy_clk
		m0_ddr3_memory_pll_sharing_pll_addr_cmd_clk                 : out   std_logic;                                        --                                     .pll_addr_cmd_clk
		m0_ddr3_memory_pll_sharing_pll_avl_clk                      : out   std_logic;                                        --                                     .pll_avl_clk
		m0_ddr3_memory_pll_sharing_pll_config_clk                   : out   std_logic;                                        --                                     .pll_config_clk
		m0_ddr3_memory_status_local_init_done                       : out   std_logic;                                        --                m0_ddr3_memory_status.local_init_done
		m0_ddr3_memory_status_local_cal_success                     : out   std_logic;                                        --                                     .local_cal_success
		m0_ddr3_memory_status_local_cal_fail                        : out   std_logic;                                        --                                     .local_cal_fail
		m0_ddr3_oct_rdn                                             : in    std_logic                     := '0';             --                          m0_ddr3_oct.rdn
		m0_ddr3_oct_rup                                             : in    std_logic                     := '0';             --                                     .rup
		rst_reset_n                                                 : in    std_logic                     := '0';             --                                  rst.reset_n
		rst_controller_conduit_reset_input_t_reset_input_signal     : in    std_logic                     := '0';             --   rst_controller_conduit_reset_input.t_reset_input_signal
		rst_controller_conduit_simucam_reset_t_simucam_reset_signal : out   std_logic;                                        -- rst_controller_conduit_simucam_reset.t_simucam_reset_signal
		sd_card_wp_n_io_export                                      : in    std_logic                     := '0';             --                      sd_card_wp_n_io.export
		slide_sw_export                                             : in    std_logic_vector(3 downto 0)  := (others => '0'); --                             slide_sw.export
		temp_scl_export                                             : out   std_logic;                                        --                             temp_scl.export
		temp_sda_export                                             : inout std_logic                     := '0';             --                             temp_sda.export
		timer_1ms_external_port_export                              : out   std_logic;                                        --              timer_1ms_external_port.export
		timer_1us_external_port_export                              : out   std_logic;                                        --              timer_1us_external_port.export
		tristate_conduit_tcm_address_out                            : out   std_logic_vector(25 downto 0);                    --                     tristate_conduit.tcm_address_out
		tristate_conduit_tcm_read_n_out                             : out   std_logic_vector(0 downto 0);                     --                                     .tcm_read_n_out
		tristate_conduit_tcm_write_n_out                            : out   std_logic_vector(0 downto 0);                     --                                     .tcm_write_n_out
		tristate_conduit_tcm_data_out                               : inout std_logic_vector(15 downto 0) := (others => '0'); --                                     .tcm_data_out
		tristate_conduit_tcm_chipselect_n_out                       : out   std_logic_vector(0 downto 0)                      --                                     .tcm_chipselect_n_out
	);
end entity MebX_Qsys_Project;

architecture rtl of MebX_Qsys_Project is
	component mfil_memory_filler_top is
		port (
			clock_sink_clk_i                  : in  std_logic                      := 'X';             -- clk
			reset_sink_reset_i                : in  std_logic                      := 'X';             -- reset
			avalon_slave_config_address_i     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avalon_slave_config_byteenable_i  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			avalon_slave_config_write_i       : in  std_logic                      := 'X';             -- write
			avalon_slave_config_writedata_i   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avalon_slave_config_read_i        : in  std_logic                      := 'X';             -- read
			avalon_slave_config_readdata_o    : out std_logic_vector(31 downto 0);                     -- readdata
			avalon_slave_config_waitrequest_o : out std_logic;                                         -- waitrequest
			avalon_master_data_waitrequest_i  : in  std_logic                      := 'X';             -- waitrequest
			avalon_master_data_address_o      : out std_logic_vector(63 downto 0);                     -- address
			avalon_master_data_write_o        : out std_logic;                                         -- write
			avalon_master_data_writedata_o    : out std_logic_vector(255 downto 0)                     -- writedata
		);
	end component mfil_memory_filler_top;

	component MebX_Qsys_Project_board_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_board_led;

	component MebX_Qsys_Project_button is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component MebX_Qsys_Project_button;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(11 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component MebX_Qsys_Project_csense_adc_fo is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_csense_adc_fo;

	component MebX_Qsys_Project_csense_cs_n is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_csense_cs_n;

	component MebX_Qsys_Project_csense_sdo is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_csense_sdo;

	component altera_address_span_extender is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			avs_s0_address       : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                     := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                     := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_readdatavalid : out std_logic;                                        -- readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_burstcount    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_m0_read          : out std_logic;                                        -- read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                        -- write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_m0_burstcount    : out std_logic_vector(7 downto 0);                     -- burstcount
			avs_cntl_read        : in  std_logic                     := 'X';             -- read
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);                    -- readdata
			avs_cntl_write       : in  std_logic                     := 'X';             -- write
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- address
		);
	end component altera_address_span_extender;

	component MebX_Qsys_Project_ext_flash is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(25 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component MebX_Qsys_Project_ext_flash;

	component MebX_Qsys_Project_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_jtag_uart;

	component MebX_Qsys_Project_m0_ddr3_i2c_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_m0_ddr3_i2c_sda;

	component MebX_Qsys_Project_m0_ddr3_memory is
		port (
			pll_ref_clk               : in    std_logic                      := 'X';             -- clk
			global_reset_n            : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n              : in    std_logic                      := 'X';             -- reset_n
			afi_clk                   : out   std_logic;                                         -- clk
			afi_half_clk              : out   std_logic;                                         -- clk
			afi_reset_n               : out   std_logic;                                         -- reset_n
			afi_reset_export_n        : out   std_logic;                                         -- reset_n
			mem_a                     : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba                    : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                    : out   std_logic_vector(0 downto 0);                      -- mem_ck
			mem_ck_n                  : out   std_logic_vector(0 downto 0);                      -- mem_ck_n
			mem_cke                   : out   std_logic_vector(0 downto 0);                      -- mem_cke
			mem_cs_n                  : out   std_logic_vector(0 downto 0);                      -- mem_cs_n
			mem_dm                    : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n                 : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n                 : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n                  : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_reset_n               : out   std_logic;                                         -- mem_reset_n
			mem_dq                    : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                   : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                 : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                   : out   std_logic_vector(0 downto 0);                      -- mem_odt
			avl_ready                 : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin            : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr                  : in    std_logic_vector(24 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid           : out   std_logic;                                         -- readdatavalid
			avl_rdata                 : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata                 : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be                    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req              : in    std_logic                      := 'X';             -- read
			avl_write_req             : in    std_logic                      := 'X';             -- write
			avl_size                  : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			local_init_done           : out   std_logic;                                         -- local_init_done
			local_cal_success         : out   std_logic;                                         -- local_cal_success
			local_cal_fail            : out   std_logic;                                         -- local_cal_fail
			oct_rdn                   : in    std_logic                      := 'X';             -- rdn
			oct_rup                   : in    std_logic                      := 'X';             -- rup
			pll_mem_clk               : out   std_logic;                                         -- pll_mem_clk
			pll_write_clk             : out   std_logic;                                         -- pll_write_clk
			pll_locked                : out   std_logic;                                         -- pll_locked
			pll_write_clk_pre_phy_clk : out   std_logic;                                         -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          : out   std_logic;                                         -- pll_addr_cmd_clk
			pll_avl_clk               : out   std_logic;                                         -- pll_avl_clk
			pll_config_clk            : out   std_logic                                          -- pll_config_clk
		);
	end component MebX_Qsys_Project_m0_ddr3_memory;

	component MebX_Qsys_Project_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(31 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component MebX_Qsys_Project_nios2_gen2_0;

	component MebX_Qsys_Project_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component MebX_Qsys_Project_onchip_memory;

	component rst_controller_top is
		port (
			clock_sink_clk                          : in  std_logic                     := 'X';             -- clk
			reset_sink_reset                        : in  std_logic                     := 'X';             -- reset
			reset_source_rs232_reset                : out std_logic;                                        -- reset
			avalon_slave_rst_controller_address     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avalon_slave_rst_controller_write       : in  std_logic                     := 'X';             -- write
			avalon_slave_rst_controller_read        : in  std_logic                     := 'X';             -- read
			avalon_slave_rst_controller_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_rst_controller_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_rst_controller_waitrequest : out std_logic;                                        -- waitrequest
			simucam_reset_signal                    : out std_logic;                                        -- t_simucam_reset_signal
			reset_input_signal                      : in  std_logic                     := 'X'              -- t_reset_input_signal
		);
	end component rst_controller_top;

	component MebX_Qsys_Project_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component MebX_Qsys_Project_sysid_qsys;

	component MebX_Qsys_Project_timer_1ms is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1ms;

	component MebX_Qsys_Project_timer_1us is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1us;

	component MebX_Qsys_Project_tristate_conduit_bridge_0 is
		port (
			clk                      : in    std_logic                     := 'X';             -- clk
			reset                    : in    std_logic                     := 'X';             -- reset
			request                  : in    std_logic                     := 'X';             -- request
			grant                    : out   std_logic;                                        -- grant
			tcs_tcm_address_out      : in    std_logic_vector(25 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out         : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen       : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in          : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out          : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tcm_read_n_out           : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component MebX_Qsys_Project_tristate_conduit_bridge_0;

	component MebX_Qsys_Project_mm_interconnect_0 is
		port (
			clk_100_clk_clk                                                 : in  std_logic                      := 'X';             -- clk
			m0_ddr3_memory_afi_clk_clk                                      : in  std_logic                      := 'X';             -- clk
			m0_ddr3_memory_avl_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			m0_ddr3_memory_soft_reset_reset_bridge_in_reset_reset           : in  std_logic                      := 'X';             -- reset
			Memory_Filler_reset_sink_reset_bridge_in_reset_reset            : in  std_logic                      := 'X';             -- reset
			ddr2_address_span_extender_expanded_master_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			ddr2_address_span_extender_expanded_master_waitrequest          : out std_logic;                                         -- waitrequest
			ddr2_address_span_extender_expanded_master_burstcount           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			ddr2_address_span_extender_expanded_master_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			ddr2_address_span_extender_expanded_master_read                 : in  std_logic                      := 'X';             -- read
			ddr2_address_span_extender_expanded_master_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			ddr2_address_span_extender_expanded_master_readdatavalid        : out std_logic;                                         -- readdatavalid
			ddr2_address_span_extender_expanded_master_write                : in  std_logic                      := 'X';             -- write
			ddr2_address_span_extender_expanded_master_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			Memory_Filler_avalon_master_data_address                        : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			Memory_Filler_avalon_master_data_waitrequest                    : out std_logic;                                         -- waitrequest
			Memory_Filler_avalon_master_data_write                          : in  std_logic                      := 'X';             -- write
			Memory_Filler_avalon_master_data_writedata                      : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			m0_ddr3_memory_avl_address                                      : out std_logic_vector(24 downto 0);                     -- address
			m0_ddr3_memory_avl_write                                        : out std_logic;                                         -- write
			m0_ddr3_memory_avl_read                                         : out std_logic;                                         -- read
			m0_ddr3_memory_avl_readdata                                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m0_ddr3_memory_avl_writedata                                    : out std_logic_vector(255 downto 0);                    -- writedata
			m0_ddr3_memory_avl_beginbursttransfer                           : out std_logic;                                         -- beginbursttransfer
			m0_ddr3_memory_avl_burstcount                                   : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_ddr3_memory_avl_byteenable                                   : out std_logic_vector(31 downto 0);                     -- byteenable
			m0_ddr3_memory_avl_readdatavalid                                : in  std_logic                      := 'X';             -- readdatavalid
			m0_ddr3_memory_avl_waitrequest                                  : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_0;

	component MebX_Qsys_Project_mm_interconnect_1 is
		port (
			clk_100_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			ext_flash_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                          : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_burstcount              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			nios2_gen2_0_instruction_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			clock_bridge_afi_50_s0_address                          : out std_logic_vector(11 downto 0);                    -- address
			clock_bridge_afi_50_s0_write                            : out std_logic;                                        -- write
			clock_bridge_afi_50_s0_read                             : out std_logic;                                        -- read
			clock_bridge_afi_50_s0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clock_bridge_afi_50_s0_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			clock_bridge_afi_50_s0_burstcount                       : out std_logic_vector(0 downto 0);                     -- burstcount
			clock_bridge_afi_50_s0_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			clock_bridge_afi_50_s0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			clock_bridge_afi_50_s0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			clock_bridge_afi_50_s0_debugaccess                      : out std_logic;                                        -- debugaccess
			ddr2_address_span_extender_cntl_write                   : out std_logic;                                        -- write
			ddr2_address_span_extender_cntl_read                    : out std_logic;                                        -- read
			ddr2_address_span_extender_cntl_readdata                : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			ddr2_address_span_extender_cntl_writedata               : out std_logic_vector(63 downto 0);                    -- writedata
			ddr2_address_span_extender_cntl_byteenable              : out std_logic_vector(7 downto 0);                     -- byteenable
			ddr2_address_span_extender_windowed_slave_address       : out std_logic_vector(28 downto 0);                    -- address
			ddr2_address_span_extender_windowed_slave_write         : out std_logic;                                        -- write
			ddr2_address_span_extender_windowed_slave_read          : out std_logic;                                        -- read
			ddr2_address_span_extender_windowed_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ddr2_address_span_extender_windowed_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			ddr2_address_span_extender_windowed_slave_burstcount    : out std_logic_vector(7 downto 0);                     -- burstcount
			ddr2_address_span_extender_windowed_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			ext_flash_uas_address                                   : out std_logic_vector(25 downto 0);                    -- address
			ext_flash_uas_write                                     : out std_logic;                                        -- write
			ext_flash_uas_read                                      : out std_logic;                                        -- read
			ext_flash_uas_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			ext_flash_uas_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			ext_flash_uas_burstcount                                : out std_logic_vector(1 downto 0);                     -- burstcount
			ext_flash_uas_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			ext_flash_uas_readdatavalid                             : in  std_logic                     := 'X';             -- readdatavalid
			ext_flash_uas_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			ext_flash_uas_lock                                      : out std_logic;                                        -- lock
			ext_flash_uas_debugaccess                               : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                  : out std_logic;                                        -- chipselect
			Memory_Filler_avalon_slave_config_address               : out std_logic_vector(7 downto 0);                     -- address
			Memory_Filler_avalon_slave_config_write                 : out std_logic;                                        -- write
			Memory_Filler_avalon_slave_config_read                  : out std_logic;                                        -- read
			Memory_Filler_avalon_slave_config_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Memory_Filler_avalon_slave_config_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			Memory_Filler_avalon_slave_config_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			Memory_Filler_avalon_slave_config_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_address                    : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                      : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                       : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                                : out std_logic_vector(17 downto 0);                    -- address
			onchip_memory_s1_write                                  : out std_logic;                                        -- write
			onchip_memory_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                                  : out std_logic;                                        -- clken
			sysid_qsys_control_slave_address                        : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component MebX_Qsys_Project_mm_interconnect_1;

	component MebX_Qsys_Project_mm_interconnect_2 is
		port (
			clk_50_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			clock_bridge_afi_50_m0_address                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_bridge_afi_50_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			clock_bridge_afi_50_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_bridge_afi_50_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_bridge_afi_50_m0_read                              : in  std_logic                     := 'X';             -- read
			clock_bridge_afi_50_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			clock_bridge_afi_50_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			clock_bridge_afi_50_m0_write                             : in  std_logic                     := 'X';             -- write
			clock_bridge_afi_50_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_bridge_afi_50_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			board_led_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			board_led_s1_write                                       : out std_logic;                                        -- write
			board_led_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			board_led_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			board_led_s1_chipselect                                  : out std_logic;                                        -- chipselect
			button_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			button_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_adc_fo_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			csense_adc_fo_s1_write                                   : out std_logic;                                        -- write
			csense_adc_fo_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_adc_fo_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			csense_adc_fo_s1_chipselect                              : out std_logic;                                        -- chipselect
			csense_cs_n_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			csense_cs_n_s1_write                                     : out std_logic;                                        -- write
			csense_cs_n_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_cs_n_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			csense_cs_n_s1_chipselect                                : out std_logic;                                        -- chipselect
			csense_sck_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			csense_sck_s1_write                                      : out std_logic;                                        -- write
			csense_sck_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sck_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sck_s1_chipselect                                 : out std_logic;                                        -- chipselect
			csense_sdi_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			csense_sdi_s1_write                                      : out std_logic;                                        -- write
			csense_sdi_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sdi_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sdi_s1_chipselect                                 : out std_logic;                                        -- chipselect
			csense_sdo_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			csense_sdo_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_ddr3_i2c_scl_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			m0_ddr3_i2c_scl_s1_write                                 : out std_logic;                                        -- write
			m0_ddr3_i2c_scl_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_ddr3_i2c_scl_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			m0_ddr3_i2c_scl_s1_chipselect                            : out std_logic;                                        -- chipselect
			m0_ddr3_i2c_sda_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			m0_ddr3_i2c_sda_s1_write                                 : out std_logic;                                        -- write
			m0_ddr3_i2c_sda_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_ddr3_i2c_sda_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			m0_ddr3_i2c_sda_s1_chipselect                            : out std_logic;                                        -- chipselect
			rst_controller_avalon_rst_controller_slave_address       : out std_logic_vector(3 downto 0);                     -- address
			rst_controller_avalon_rst_controller_slave_write         : out std_logic;                                        -- write
			rst_controller_avalon_rst_controller_slave_read          : out std_logic;                                        -- read
			rst_controller_avalon_rst_controller_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rst_controller_avalon_rst_controller_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			rst_controller_avalon_rst_controller_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			sd_card_wp_n_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			sd_card_wp_n_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			slide_sw_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			slide_sw_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_scl_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			temp_scl_s1_write                                        : out std_logic;                                        -- write
			temp_scl_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_scl_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			temp_scl_s1_chipselect                                   : out std_logic;                                        -- chipselect
			temp_sda_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			temp_sda_s1_write                                        : out std_logic;                                        -- write
			temp_sda_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_sda_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			temp_sda_s1_chipselect                                   : out std_logic;                                        -- chipselect
			timer_1ms_s1_address                                     : out std_logic_vector(2 downto 0);                     -- address
			timer_1ms_s1_write                                       : out std_logic;                                        -- write
			timer_1ms_s1_readdata                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1ms_s1_writedata                                   : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1ms_s1_chipselect                                  : out std_logic;                                        -- chipselect
			timer_1us_s1_address                                     : out std_logic_vector(2 downto 0);                     -- address
			timer_1us_s1_write                                       : out std_logic;                                        -- write
			timer_1us_s1_readdata                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1us_s1_writedata                                   : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1us_s1_chipselect                                  : out std_logic                                         -- chipselect
		);
	end component MebX_Qsys_Project_mm_interconnect_2;

	component MebX_Qsys_Project_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component MebX_Qsys_Project_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component mebx_qsys_project_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_001;

	component mebx_qsys_project_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_002;

	component mebx_qsys_project_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_003;

	signal m0_ddr3_memory_afi_clk_clk                                                : std_logic;                      -- m0_ddr3_memory:afi_clk -> [mm_interconnect_0:m0_ddr3_memory_afi_clk_clk, rst_controller_005:clk]
	signal m0_ddr3_memory_afi_half_clk_clk                                           : std_logic;                      -- m0_ddr3_memory:afi_half_clk -> [Memory_Filler:clock_sink_clk_i, clock_bridge_afi_50:s0_clk, ddr2_address_span_extender:clk, ext_flash:clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:clk_100_clk_clk, mm_interconnect_1:clk_100_clk_clk, nios2_gen2_0:clk, onchip_memory:clk, rst_controller_001:clk, rst_controller_003:clk, rst_controller_004:clk, sysid_qsys:clock, tristate_conduit_bridge_0:clk]
	signal ext_flash_tcm_data_outen                                                  : std_logic;                      -- ext_flash:tcm_data_outen -> tristate_conduit_bridge_0:tcs_tcm_data_outen
	signal ext_flash_tcm_request                                                     : std_logic;                      -- ext_flash:tcm_request -> tristate_conduit_bridge_0:request
	signal ext_flash_tcm_write_n_out                                                 : std_logic;                      -- ext_flash:tcm_write_n_out -> tristate_conduit_bridge_0:tcs_tcm_write_n_out
	signal ext_flash_tcm_read_n_out                                                  : std_logic;                      -- ext_flash:tcm_read_n_out -> tristate_conduit_bridge_0:tcs_tcm_read_n_out
	signal ext_flash_tcm_grant                                                       : std_logic;                      -- tristate_conduit_bridge_0:grant -> ext_flash:tcm_grant
	signal ext_flash_tcm_chipselect_n_out                                            : std_logic;                      -- ext_flash:tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_tcm_chipselect_n_out
	signal ext_flash_tcm_address_out                                                 : std_logic_vector(25 downto 0);  -- ext_flash:tcm_address_out -> tristate_conduit_bridge_0:tcs_tcm_address_out
	signal ext_flash_tcm_data_out                                                    : std_logic_vector(15 downto 0);  -- ext_flash:tcm_data_out -> tristate_conduit_bridge_0:tcs_tcm_data_out
	signal ext_flash_tcm_data_in                                                     : std_logic_vector(15 downto 0);  -- tristate_conduit_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	signal memory_filler_avalon_master_data_waitrequest                              : std_logic;                      -- mm_interconnect_0:Memory_Filler_avalon_master_data_waitrequest -> Memory_Filler:avalon_master_data_waitrequest_i
	signal memory_filler_avalon_master_data_address                                  : std_logic_vector(63 downto 0);  -- Memory_Filler:avalon_master_data_address_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_address
	signal memory_filler_avalon_master_data_write                                    : std_logic;                      -- Memory_Filler:avalon_master_data_write_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_write
	signal memory_filler_avalon_master_data_writedata                                : std_logic_vector(255 downto 0); -- Memory_Filler:avalon_master_data_writedata_o -> mm_interconnect_0:Memory_Filler_avalon_master_data_writedata
	signal ddr2_address_span_extender_expanded_master_waitrequest                    : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_waitrequest -> ddr2_address_span_extender:avm_m0_waitrequest
	signal ddr2_address_span_extender_expanded_master_readdata                       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdata -> ddr2_address_span_extender:avm_m0_readdata
	signal ddr2_address_span_extender_expanded_master_address                        : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_address -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_address
	signal ddr2_address_span_extender_expanded_master_read                           : std_logic;                      -- ddr2_address_span_extender:avm_m0_read -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_read
	signal ddr2_address_span_extender_expanded_master_byteenable                     : std_logic_vector(3 downto 0);   -- ddr2_address_span_extender:avm_m0_byteenable -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_byteenable
	signal ddr2_address_span_extender_expanded_master_readdatavalid                  : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdatavalid -> ddr2_address_span_extender:avm_m0_readdatavalid
	signal ddr2_address_span_extender_expanded_master_write                          : std_logic;                      -- ddr2_address_span_extender:avm_m0_write -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_write
	signal ddr2_address_span_extender_expanded_master_writedata                      : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_writedata -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_writedata
	signal ddr2_address_span_extender_expanded_master_burstcount                     : std_logic_vector(7 downto 0);   -- ddr2_address_span_extender:avm_m0_burstcount -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_burstcount
	signal mm_interconnect_0_m0_ddr3_memory_avl_beginbursttransfer                   : std_logic;                      -- mm_interconnect_0:m0_ddr3_memory_avl_beginbursttransfer -> m0_ddr3_memory:avl_burstbegin
	signal mm_interconnect_0_m0_ddr3_memory_avl_readdata                             : std_logic_vector(255 downto 0); -- m0_ddr3_memory:avl_rdata -> mm_interconnect_0:m0_ddr3_memory_avl_readdata
	signal m0_ddr3_memory_avl_waitrequest                                            : std_logic;                      -- m0_ddr3_memory:avl_ready -> m0_ddr3_memory_avl_waitrequest:in
	signal mm_interconnect_0_m0_ddr3_memory_avl_address                              : std_logic_vector(24 downto 0);  -- mm_interconnect_0:m0_ddr3_memory_avl_address -> m0_ddr3_memory:avl_addr
	signal mm_interconnect_0_m0_ddr3_memory_avl_read                                 : std_logic;                      -- mm_interconnect_0:m0_ddr3_memory_avl_read -> m0_ddr3_memory:avl_read_req
	signal mm_interconnect_0_m0_ddr3_memory_avl_byteenable                           : std_logic_vector(31 downto 0);  -- mm_interconnect_0:m0_ddr3_memory_avl_byteenable -> m0_ddr3_memory:avl_be
	signal mm_interconnect_0_m0_ddr3_memory_avl_readdatavalid                        : std_logic;                      -- m0_ddr3_memory:avl_rdata_valid -> mm_interconnect_0:m0_ddr3_memory_avl_readdatavalid
	signal mm_interconnect_0_m0_ddr3_memory_avl_write                                : std_logic;                      -- mm_interconnect_0:m0_ddr3_memory_avl_write -> m0_ddr3_memory:avl_write_req
	signal mm_interconnect_0_m0_ddr3_memory_avl_writedata                            : std_logic_vector(255 downto 0); -- mm_interconnect_0:m0_ddr3_memory_avl_writedata -> m0_ddr3_memory:avl_wdata
	signal mm_interconnect_0_m0_ddr3_memory_avl_burstcount                           : std_logic_vector(3 downto 0);   -- mm_interconnect_0:m0_ddr3_memory_avl_burstcount -> m0_ddr3_memory:avl_size
	signal nios2_gen2_0_data_master_readdata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                      : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                      : std_logic;                      -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                          : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                       : std_logic_vector(3 downto 0);   -- nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                             : std_logic;                      -- nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                            : std_logic;                      -- nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                        : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                               : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                   : std_logic_vector(31 downto 0);  -- nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                      : std_logic;                      -- nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                             : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal nios2_gen2_0_instruction_master_burstcount                                : std_logic_vector(3 downto 0);   -- nios2_gen2_0:i_burstcount -> mm_interconnect_1:nios2_gen2_0_instruction_master_burstcount
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect                  : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata                    : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest                 : std_logic;                      -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address                     : std_logic_vector(0 downto 0);   -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read                        : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write                       : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_memory_filler_avalon_slave_config_readdata              : std_logic_vector(31 downto 0);  -- Memory_Filler:avalon_slave_config_readdata_o -> mm_interconnect_1:Memory_Filler_avalon_slave_config_readdata
	signal mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest           : std_logic;                      -- Memory_Filler:avalon_slave_config_waitrequest_o -> mm_interconnect_1:Memory_Filler_avalon_slave_config_waitrequest
	signal mm_interconnect_1_memory_filler_avalon_slave_config_address               : std_logic_vector(7 downto 0);   -- mm_interconnect_1:Memory_Filler_avalon_slave_config_address -> Memory_Filler:avalon_slave_config_address_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_read                  : std_logic;                      -- mm_interconnect_1:Memory_Filler_avalon_slave_config_read -> Memory_Filler:avalon_slave_config_read_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_byteenable            : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Memory_Filler_avalon_slave_config_byteenable -> Memory_Filler:avalon_slave_config_byteenable_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_write                 : std_logic;                      -- mm_interconnect_1:Memory_Filler_avalon_slave_config_write -> Memory_Filler:avalon_slave_config_write_i
	signal mm_interconnect_1_memory_filler_avalon_slave_config_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Memory_Filler_avalon_slave_config_writedata -> Memory_Filler:avalon_slave_config_writedata_i
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_readdata                : std_logic_vector(63 downto 0);  -- ddr2_address_span_extender:avs_cntl_readdata -> mm_interconnect_1:ddr2_address_span_extender_cntl_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_read                    : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_read -> ddr2_address_span_extender:avs_cntl_read
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable              : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_cntl_byteenable -> ddr2_address_span_extender:avs_cntl_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_write                   : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_write -> ddr2_address_span_extender:avs_cntl_write
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_writedata               : std_logic_vector(63 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_cntl_writedata -> ddr2_address_span_extender:avs_cntl_writedata
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata                       : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address                        : std_logic_vector(0 downto 0);   -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata                   : std_logic_vector(31 downto 0);  -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest                : std_logic;                      -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess                : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address                    : std_logic_vector(8 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read                       : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable                 : std_logic_vector(3 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write                      : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata                  : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdata                         : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:s0_readdata -> mm_interconnect_1:clock_bridge_afi_50_s0_readdata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest                      : std_logic;                      -- clock_bridge_afi_50:s0_waitrequest -> mm_interconnect_1:clock_bridge_afi_50_s0_waitrequest
	signal mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess                      : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_debugaccess -> clock_bridge_afi_50:s0_debugaccess
	signal mm_interconnect_1_clock_bridge_afi_50_s0_address                          : std_logic_vector(11 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_address -> clock_bridge_afi_50:s0_address
	signal mm_interconnect_1_clock_bridge_afi_50_s0_read                             : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_read -> clock_bridge_afi_50:s0_read
	signal mm_interconnect_1_clock_bridge_afi_50_s0_byteenable                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_byteenable -> clock_bridge_afi_50:s0_byteenable
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid                    : std_logic;                      -- clock_bridge_afi_50:s0_readdatavalid -> mm_interconnect_1:clock_bridge_afi_50_s0_readdatavalid
	signal mm_interconnect_1_clock_bridge_afi_50_s0_write                            : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_write -> clock_bridge_afi_50:s0_write
	signal mm_interconnect_1_clock_bridge_afi_50_s0_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_writedata -> clock_bridge_afi_50:s0_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_burstcount                       : std_logic_vector(0 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_burstcount -> clock_bridge_afi_50:s0_burstcount
	signal mm_interconnect_1_onchip_memory_s1_chipselect                             : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_1_onchip_memory_s1_readdata                               : std_logic_vector(31 downto 0);  -- onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	signal mm_interconnect_1_onchip_memory_s1_address                                : std_logic_vector(17 downto 0);  -- mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_1_onchip_memory_s1_byteenable                             : std_logic_vector(3 downto 0);   -- mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_1_onchip_memory_s1_write                                  : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_1_onchip_memory_s1_writedata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_1_onchip_memory_s1_clken                                  : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_1_ext_flash_uas_readdata                                  : std_logic_vector(15 downto 0);  -- ext_flash:uas_readdata -> mm_interconnect_1:ext_flash_uas_readdata
	signal mm_interconnect_1_ext_flash_uas_waitrequest                               : std_logic;                      -- ext_flash:uas_waitrequest -> mm_interconnect_1:ext_flash_uas_waitrequest
	signal mm_interconnect_1_ext_flash_uas_debugaccess                               : std_logic;                      -- mm_interconnect_1:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	signal mm_interconnect_1_ext_flash_uas_address                                   : std_logic_vector(25 downto 0);  -- mm_interconnect_1:ext_flash_uas_address -> ext_flash:uas_address
	signal mm_interconnect_1_ext_flash_uas_read                                      : std_logic;                      -- mm_interconnect_1:ext_flash_uas_read -> ext_flash:uas_read
	signal mm_interconnect_1_ext_flash_uas_byteenable                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	signal mm_interconnect_1_ext_flash_uas_readdatavalid                             : std_logic;                      -- ext_flash:uas_readdatavalid -> mm_interconnect_1:ext_flash_uas_readdatavalid
	signal mm_interconnect_1_ext_flash_uas_lock                                      : std_logic;                      -- mm_interconnect_1:ext_flash_uas_lock -> ext_flash:uas_lock
	signal mm_interconnect_1_ext_flash_uas_write                                     : std_logic;                      -- mm_interconnect_1:ext_flash_uas_write -> ext_flash:uas_write
	signal mm_interconnect_1_ext_flash_uas_writedata                                 : std_logic_vector(15 downto 0);  -- mm_interconnect_1:ext_flash_uas_writedata -> ext_flash:uas_writedata
	signal mm_interconnect_1_ext_flash_uas_burstcount                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata      : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avs_s0_readdata -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest   : std_logic;                      -- ddr2_address_span_extender:avs_s0_waitrequest -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_waitrequest
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address       : std_logic_vector(28 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_address -> ddr2_address_span_extender:avs_s0_address
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read          : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_read -> ddr2_address_span_extender:avs_s0_read
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable    : std_logic_vector(3 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_byteenable -> ddr2_address_span_extender:avs_s0_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid : std_logic;                      -- ddr2_address_span_extender:avs_s0_readdatavalid -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdatavalid
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write         : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_write -> ddr2_address_span_extender:avs_s0_write
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_writedata -> ddr2_address_span_extender:avs_s0_writedata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount    : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_burstcount -> ddr2_address_span_extender:avs_s0_burstcount
	signal clock_bridge_afi_50_m0_waitrequest                                        : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_waitrequest -> clock_bridge_afi_50:m0_waitrequest
	signal clock_bridge_afi_50_m0_readdata                                           : std_logic_vector(31 downto 0);  -- mm_interconnect_2:clock_bridge_afi_50_m0_readdata -> clock_bridge_afi_50:m0_readdata
	signal clock_bridge_afi_50_m0_debugaccess                                        : std_logic;                      -- clock_bridge_afi_50:m0_debugaccess -> mm_interconnect_2:clock_bridge_afi_50_m0_debugaccess
	signal clock_bridge_afi_50_m0_address                                            : std_logic_vector(11 downto 0);  -- clock_bridge_afi_50:m0_address -> mm_interconnect_2:clock_bridge_afi_50_m0_address
	signal clock_bridge_afi_50_m0_read                                               : std_logic;                      -- clock_bridge_afi_50:m0_read -> mm_interconnect_2:clock_bridge_afi_50_m0_read
	signal clock_bridge_afi_50_m0_byteenable                                         : std_logic_vector(3 downto 0);   -- clock_bridge_afi_50:m0_byteenable -> mm_interconnect_2:clock_bridge_afi_50_m0_byteenable
	signal clock_bridge_afi_50_m0_readdatavalid                                      : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_readdatavalid -> clock_bridge_afi_50:m0_readdatavalid
	signal clock_bridge_afi_50_m0_writedata                                          : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:m0_writedata -> mm_interconnect_2:clock_bridge_afi_50_m0_writedata
	signal clock_bridge_afi_50_m0_write                                              : std_logic;                      -- clock_bridge_afi_50:m0_write -> mm_interconnect_2:clock_bridge_afi_50_m0_write
	signal clock_bridge_afi_50_m0_burstcount                                         : std_logic_vector(0 downto 0);   -- clock_bridge_afi_50:m0_burstcount -> mm_interconnect_2:clock_bridge_afi_50_m0_burstcount
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata     : std_logic_vector(31 downto 0);  -- rst_controller:avalon_slave_rst_controller_readdata -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_readdata
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest  : std_logic;                      -- rst_controller:avalon_slave_rst_controller_waitrequest -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_waitrequest
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address      : std_logic_vector(3 downto 0);   -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_address -> rst_controller:avalon_slave_rst_controller_address
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read         : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_read -> rst_controller:avalon_slave_rst_controller_read
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write        : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_write -> rst_controller:avalon_slave_rst_controller_write
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_writedata -> rst_controller:avalon_slave_rst_controller_writedata
	signal mm_interconnect_2_timer_1ms_s1_chipselect                                 : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_chipselect -> timer_1ms:chipselect
	signal mm_interconnect_2_timer_1ms_s1_readdata                                   : std_logic_vector(15 downto 0);  -- timer_1ms:readdata -> mm_interconnect_2:timer_1ms_s1_readdata
	signal mm_interconnect_2_timer_1ms_s1_address                                    : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1ms_s1_address -> timer_1ms:address
	signal mm_interconnect_2_timer_1ms_s1_write                                      : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_write -> mm_interconnect_2_timer_1ms_s1_write:in
	signal mm_interconnect_2_timer_1ms_s1_writedata                                  : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1ms_s1_writedata -> timer_1ms:writedata
	signal mm_interconnect_2_timer_1us_s1_chipselect                                 : std_logic;                      -- mm_interconnect_2:timer_1us_s1_chipselect -> timer_1us:chipselect
	signal mm_interconnect_2_timer_1us_s1_readdata                                   : std_logic_vector(15 downto 0);  -- timer_1us:readdata -> mm_interconnect_2:timer_1us_s1_readdata
	signal mm_interconnect_2_timer_1us_s1_address                                    : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1us_s1_address -> timer_1us:address
	signal mm_interconnect_2_timer_1us_s1_write                                      : std_logic;                      -- mm_interconnect_2:timer_1us_s1_write -> mm_interconnect_2_timer_1us_s1_write:in
	signal mm_interconnect_2_timer_1us_s1_writedata                                  : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1us_s1_writedata -> timer_1us:writedata
	signal mm_interconnect_2_sd_card_wp_n_s1_readdata                                : std_logic_vector(31 downto 0);  -- sd_card_wp_n:readdata -> mm_interconnect_2:sd_card_wp_n_s1_readdata
	signal mm_interconnect_2_sd_card_wp_n_s1_address                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_2:sd_card_wp_n_s1_address -> sd_card_wp_n:address
	signal mm_interconnect_2_temp_scl_s1_chipselect                                  : std_logic;                      -- mm_interconnect_2:temp_scl_s1_chipselect -> temp_scl:chipselect
	signal mm_interconnect_2_temp_scl_s1_readdata                                    : std_logic_vector(31 downto 0);  -- temp_scl:readdata -> mm_interconnect_2:temp_scl_s1_readdata
	signal mm_interconnect_2_temp_scl_s1_address                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_scl_s1_address -> temp_scl:address
	signal mm_interconnect_2_temp_scl_s1_write                                       : std_logic;                      -- mm_interconnect_2:temp_scl_s1_write -> mm_interconnect_2_temp_scl_s1_write:in
	signal mm_interconnect_2_temp_scl_s1_writedata                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_scl_s1_writedata -> temp_scl:writedata
	signal mm_interconnect_2_temp_sda_s1_chipselect                                  : std_logic;                      -- mm_interconnect_2:temp_sda_s1_chipselect -> temp_sda:chipselect
	signal mm_interconnect_2_temp_sda_s1_readdata                                    : std_logic_vector(31 downto 0);  -- temp_sda:readdata -> mm_interconnect_2:temp_sda_s1_readdata
	signal mm_interconnect_2_temp_sda_s1_address                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_sda_s1_address -> temp_sda:address
	signal mm_interconnect_2_temp_sda_s1_write                                       : std_logic;                      -- mm_interconnect_2:temp_sda_s1_write -> mm_interconnect_2_temp_sda_s1_write:in
	signal mm_interconnect_2_temp_sda_s1_writedata                                   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_sda_s1_writedata -> temp_sda:writedata
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_chipselect                           : std_logic;                      -- mm_interconnect_2:m0_ddr3_i2c_sda_s1_chipselect -> m0_ddr3_i2c_sda:chipselect
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_readdata                             : std_logic_vector(31 downto 0);  -- m0_ddr3_i2c_sda:readdata -> mm_interconnect_2:m0_ddr3_i2c_sda_s1_readdata
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_address                              : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m0_ddr3_i2c_sda_s1_address -> m0_ddr3_i2c_sda:address
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_write                                : std_logic;                      -- mm_interconnect_2:m0_ddr3_i2c_sda_s1_write -> mm_interconnect_2_m0_ddr3_i2c_sda_s1_write:in
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_writedata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m0_ddr3_i2c_sda_s1_writedata -> m0_ddr3_i2c_sda:writedata
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_chipselect                           : std_logic;                      -- mm_interconnect_2:m0_ddr3_i2c_scl_s1_chipselect -> m0_ddr3_i2c_scl:chipselect
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_readdata                             : std_logic_vector(31 downto 0);  -- m0_ddr3_i2c_scl:readdata -> mm_interconnect_2:m0_ddr3_i2c_scl_s1_readdata
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_address                              : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m0_ddr3_i2c_scl_s1_address -> m0_ddr3_i2c_scl:address
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_write                                : std_logic;                      -- mm_interconnect_2:m0_ddr3_i2c_scl_s1_write -> mm_interconnect_2_m0_ddr3_i2c_scl_s1_write:in
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_writedata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m0_ddr3_i2c_scl_s1_writedata -> m0_ddr3_i2c_scl:writedata
	signal mm_interconnect_2_csense_sdo_s1_readdata                                  : std_logic_vector(31 downto 0);  -- csense_sdo:readdata -> mm_interconnect_2:csense_sdo_s1_readdata
	signal mm_interconnect_2_csense_sdo_s1_address                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdo_s1_address -> csense_sdo:address
	signal mm_interconnect_2_csense_sdi_s1_chipselect                                : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_chipselect -> csense_sdi:chipselect
	signal mm_interconnect_2_csense_sdi_s1_readdata                                  : std_logic_vector(31 downto 0);  -- csense_sdi:readdata -> mm_interconnect_2:csense_sdi_s1_readdata
	signal mm_interconnect_2_csense_sdi_s1_address                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdi_s1_address -> csense_sdi:address
	signal mm_interconnect_2_csense_sdi_s1_write                                     : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_write -> mm_interconnect_2_csense_sdi_s1_write:in
	signal mm_interconnect_2_csense_sdi_s1_writedata                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sdi_s1_writedata -> csense_sdi:writedata
	signal mm_interconnect_2_csense_sck_s1_chipselect                                : std_logic;                      -- mm_interconnect_2:csense_sck_s1_chipselect -> csense_sck:chipselect
	signal mm_interconnect_2_csense_sck_s1_readdata                                  : std_logic_vector(31 downto 0);  -- csense_sck:readdata -> mm_interconnect_2:csense_sck_s1_readdata
	signal mm_interconnect_2_csense_sck_s1_address                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sck_s1_address -> csense_sck:address
	signal mm_interconnect_2_csense_sck_s1_write                                     : std_logic;                      -- mm_interconnect_2:csense_sck_s1_write -> mm_interconnect_2_csense_sck_s1_write:in
	signal mm_interconnect_2_csense_sck_s1_writedata                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sck_s1_writedata -> csense_sck:writedata
	signal mm_interconnect_2_csense_cs_n_s1_chipselect                               : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_chipselect -> csense_cs_n:chipselect
	signal mm_interconnect_2_csense_cs_n_s1_readdata                                 : std_logic_vector(31 downto 0);  -- csense_cs_n:readdata -> mm_interconnect_2:csense_cs_n_s1_readdata
	signal mm_interconnect_2_csense_cs_n_s1_address                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_cs_n_s1_address -> csense_cs_n:address
	signal mm_interconnect_2_csense_cs_n_s1_write                                    : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_write -> mm_interconnect_2_csense_cs_n_s1_write:in
	signal mm_interconnect_2_csense_cs_n_s1_writedata                                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_cs_n_s1_writedata -> csense_cs_n:writedata
	signal mm_interconnect_2_csense_adc_fo_s1_chipselect                             : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_chipselect -> csense_adc_fo:chipselect
	signal mm_interconnect_2_csense_adc_fo_s1_readdata                               : std_logic_vector(31 downto 0);  -- csense_adc_fo:readdata -> mm_interconnect_2:csense_adc_fo_s1_readdata
	signal mm_interconnect_2_csense_adc_fo_s1_address                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_adc_fo_s1_address -> csense_adc_fo:address
	signal mm_interconnect_2_csense_adc_fo_s1_write                                  : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_write -> mm_interconnect_2_csense_adc_fo_s1_write:in
	signal mm_interconnect_2_csense_adc_fo_s1_writedata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_adc_fo_s1_writedata -> csense_adc_fo:writedata
	signal mm_interconnect_2_button_s1_readdata                                      : std_logic_vector(31 downto 0);  -- button:readdata -> mm_interconnect_2:button_s1_readdata
	signal mm_interconnect_2_button_s1_address                                       : std_logic_vector(1 downto 0);   -- mm_interconnect_2:button_s1_address -> button:address
	signal mm_interconnect_2_slide_sw_s1_readdata                                    : std_logic_vector(31 downto 0);  -- slide_sw:readdata -> mm_interconnect_2:slide_sw_s1_readdata
	signal mm_interconnect_2_slide_sw_s1_address                                     : std_logic_vector(1 downto 0);   -- mm_interconnect_2:slide_sw_s1_address -> slide_sw:address
	signal mm_interconnect_2_board_led_s1_chipselect                                 : std_logic;                      -- mm_interconnect_2:board_led_s1_chipselect -> board_led:chipselect
	signal mm_interconnect_2_board_led_s1_readdata                                   : std_logic_vector(31 downto 0);  -- board_led:readdata -> mm_interconnect_2:board_led_s1_readdata
	signal mm_interconnect_2_board_led_s1_address                                    : std_logic_vector(1 downto 0);   -- mm_interconnect_2:board_led_s1_address -> board_led:address
	signal mm_interconnect_2_board_led_s1_write                                      : std_logic;                      -- mm_interconnect_2:board_led_s1_write -> mm_interconnect_2_board_led_s1_write:in
	signal mm_interconnect_2_board_led_s1_writedata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_2:board_led_s1_writedata -> board_led:writedata
	signal irq_mapper_receiver0_irq                                                  : std_logic;                      -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                                      : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver1_irq                                                  : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_receiver_irq                                             : std_logic_vector(0 downto 0);   -- timer_1ms:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver2_irq                                                  : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_001_receiver_irq                                         : std_logic_vector(0 downto 0);   -- timer_1us:irq -> irq_synchronizer_001:receiver_irq
	signal rst_controller_001_reset_out_reset                                        : std_logic;                      -- rst_controller_001:reset_out -> [Memory_Filler:reset_sink_reset_i, clock_bridge_afi_50:s0_reset, ddr2_address_span_extender:reset, mm_interconnect_0:Memory_Filler_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                                    : std_logic;                      -- rst_controller_001:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                                        : std_logic;                      -- rst_controller_002:reset_out -> [clock_bridge_afi_50:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_2:clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset, rst_controller:reset_sink_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                                        : std_logic;                      -- rst_controller_003:reset_out -> [ext_flash:reset_reset, mm_interconnect_1:ext_flash_reset_reset_bridge_in_reset_reset, tristate_conduit_bridge_0:reset]
	signal rst_controller_004_reset_out_reset                                        : std_logic;                      -- rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_004_reset_out_reset_req                                    : std_logic;                      -- rst_controller_004:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_005_reset_out_reset                                        : std_logic;                      -- rst_controller_005:reset_out -> [mm_interconnect_0:m0_ddr3_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:m0_ddr3_memory_soft_reset_reset_bridge_in_reset_reset]
	signal rst_reset_n_ports_inv                                                     : std_logic;                      -- rst_reset_n:inv -> [rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_003:reset_in1, rst_controller_004:reset_in0, rst_controller_005:reset_in0]
	signal mm_interconnect_0_m0_ddr3_memory_avl_inv                                  : std_logic;                      -- m0_ddr3_memory_avl_waitrequest:inv -> mm_interconnect_0:m0_ddr3_memory_avl_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv              : std_logic;                      -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv             : std_logic;                      -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_2_timer_1ms_s1_write_ports_inv                            : std_logic;                      -- mm_interconnect_2_timer_1ms_s1_write:inv -> timer_1ms:write_n
	signal mm_interconnect_2_timer_1us_s1_write_ports_inv                            : std_logic;                      -- mm_interconnect_2_timer_1us_s1_write:inv -> timer_1us:write_n
	signal mm_interconnect_2_temp_scl_s1_write_ports_inv                             : std_logic;                      -- mm_interconnect_2_temp_scl_s1_write:inv -> temp_scl:write_n
	signal mm_interconnect_2_temp_sda_s1_write_ports_inv                             : std_logic;                      -- mm_interconnect_2_temp_sda_s1_write:inv -> temp_sda:write_n
	signal mm_interconnect_2_m0_ddr3_i2c_sda_s1_write_ports_inv                      : std_logic;                      -- mm_interconnect_2_m0_ddr3_i2c_sda_s1_write:inv -> m0_ddr3_i2c_sda:write_n
	signal mm_interconnect_2_m0_ddr3_i2c_scl_s1_write_ports_inv                      : std_logic;                      -- mm_interconnect_2_m0_ddr3_i2c_scl_s1_write:inv -> m0_ddr3_i2c_scl:write_n
	signal mm_interconnect_2_csense_sdi_s1_write_ports_inv                           : std_logic;                      -- mm_interconnect_2_csense_sdi_s1_write:inv -> csense_sdi:write_n
	signal mm_interconnect_2_csense_sck_s1_write_ports_inv                           : std_logic;                      -- mm_interconnect_2_csense_sck_s1_write:inv -> csense_sck:write_n
	signal mm_interconnect_2_csense_cs_n_s1_write_ports_inv                          : std_logic;                      -- mm_interconnect_2_csense_cs_n_s1_write:inv -> csense_cs_n:write_n
	signal mm_interconnect_2_csense_adc_fo_s1_write_ports_inv                        : std_logic;                      -- mm_interconnect_2_csense_adc_fo_s1_write:inv -> csense_adc_fo:write_n
	signal mm_interconnect_2_board_led_s1_write_ports_inv                            : std_logic;                      -- mm_interconnect_2_board_led_s1_write:inv -> board_led:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                              : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [jtag_uart:rst_n, sysid_qsys:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                              : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> [board_led:reset_n, button:reset_n, csense_adc_fo:reset_n, csense_cs_n:reset_n, csense_sck:reset_n, csense_sdi:reset_n, csense_sdo:reset_n, m0_ddr3_i2c_scl:reset_n, m0_ddr3_i2c_sda:reset_n, sd_card_wp_n:reset_n, slide_sw:reset_n, temp_scl:reset_n, temp_sda:reset_n, timer_1ms:reset_n, timer_1us:reset_n]
	signal rst_controller_004_reset_out_reset_ports_inv                              : std_logic;                      -- rst_controller_004_reset_out_reset:inv -> nios2_gen2_0:reset_n

begin

	memory_filler : component mfil_memory_filler_top
		port map (
			clock_sink_clk_i                  => m0_ddr3_memory_afi_half_clk_clk,                                 --          clock_sink.clk
			reset_sink_reset_i                => rst_controller_001_reset_out_reset,                              --          reset_sink.reset
			avalon_slave_config_address_i     => mm_interconnect_1_memory_filler_avalon_slave_config_address,     -- avalon_slave_config.address
			avalon_slave_config_byteenable_i  => mm_interconnect_1_memory_filler_avalon_slave_config_byteenable,  --                    .byteenable
			avalon_slave_config_write_i       => mm_interconnect_1_memory_filler_avalon_slave_config_write,       --                    .write
			avalon_slave_config_writedata_i   => mm_interconnect_1_memory_filler_avalon_slave_config_writedata,   --                    .writedata
			avalon_slave_config_read_i        => mm_interconnect_1_memory_filler_avalon_slave_config_read,        --                    .read
			avalon_slave_config_readdata_o    => mm_interconnect_1_memory_filler_avalon_slave_config_readdata,    --                    .readdata
			avalon_slave_config_waitrequest_o => mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest, --                    .waitrequest
			avalon_master_data_waitrequest_i  => memory_filler_avalon_master_data_waitrequest,                    --  avalon_master_data.waitrequest
			avalon_master_data_address_o      => memory_filler_avalon_master_data_address,                        --                    .address
			avalon_master_data_write_o        => memory_filler_avalon_master_data_write,                          --                    .write
			avalon_master_data_writedata_o    => memory_filler_avalon_master_data_writedata                       --                    .writedata
		);

	board_led : component MebX_Qsys_Project_board_led
		port map (
			clk        => clk50_clk,                                      --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_2_board_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_board_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_board_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_board_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_board_led_s1_readdata,        --                    .readdata
			out_port   => board_led_export                                -- external_connection.export
		);

	button : component MebX_Qsys_Project_button
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_button_s1_address,          --                  s1.address
			readdata => mm_interconnect_2_button_s1_readdata,         --                    .readdata
			in_port  => button_export                                 -- external_connection.export
		);

	clock_bridge_afi_50 : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk50_clk,                                              --   m0_clk.clk
			m0_reset         => rst_controller_002_reset_out_reset,                     -- m0_reset.reset
			s0_clk           => m0_ddr3_memory_afi_half_clk_clk,                        --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                     -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_1_clock_bridge_afi_50_s0_address,       --         .address
			s0_write         => mm_interconnect_1_clock_bridge_afi_50_s0_write,         --         .write
			s0_read          => mm_interconnect_1_clock_bridge_afi_50_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => clock_bridge_afi_50_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => clock_bridge_afi_50_m0_readdata,                        --         .readdata
			m0_readdatavalid => clock_bridge_afi_50_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => clock_bridge_afi_50_m0_burstcount,                      --         .burstcount
			m0_writedata     => clock_bridge_afi_50_m0_writedata,                       --         .writedata
			m0_address       => clock_bridge_afi_50_m0_address,                         --         .address
			m0_write         => clock_bridge_afi_50_m0_write,                           --         .write
			m0_read          => clock_bridge_afi_50_m0_read,                            --         .read
			m0_byteenable    => clock_bridge_afi_50_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => clock_bridge_afi_50_m0_debugaccess                      --         .debugaccess
		);

	csense_adc_fo : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                          --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_2_csense_adc_fo_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_adc_fo_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_adc_fo_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_adc_fo_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_adc_fo_s1_readdata,        --                    .readdata
			out_port   => csense_adc_fo_export                                -- external_connection.export
		);

	csense_cs_n : component MebX_Qsys_Project_csense_cs_n
		port map (
			clk        => clk50_clk,                                        --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_2_csense_cs_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_cs_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_cs_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_cs_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_cs_n_s1_readdata,        --                    .readdata
			out_port   => csense_cs_n_export                                -- external_connection.export
		);

	csense_sck : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sck_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sck_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sck_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sck_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sck_s1_readdata,        --                    .readdata
			out_port   => csense_sck_export                                -- external_connection.export
		);

	csense_sdi : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sdi_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sdi_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sdi_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sdi_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sdi_s1_readdata,        --                    .readdata
			out_port   => csense_sdi_export                                -- external_connection.export
		);

	csense_sdo : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_csense_sdo_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_csense_sdo_s1_readdata,     --                    .readdata
			in_port  => csense_sdo_export                             -- external_connection.export
		);

	ddr2_address_span_extender : component altera_address_span_extender
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 29,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 8,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			clk                  => m0_ddr3_memory_afi_half_clk_clk,                                           --           clock.clk
			reset                => rst_controller_001_reset_out_reset,                                        --           reset.reset
			avs_s0_address       => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => ddr2_address_span_extender_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => ddr2_address_span_extender_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => ddr2_address_span_extender_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => ddr2_address_span_extender_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => ddr2_address_span_extender_expanded_master_write,                          --                .write
			avm_m0_writedata     => ddr2_address_span_extender_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => ddr2_address_span_extender_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => ddr2_address_span_extender_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => ddr2_address_span_extender_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_read        => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                    --            cntl.read
			avs_cntl_readdata    => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                --                .readdata
			avs_cntl_write       => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                   --                .write
			avs_cntl_writedata   => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,               --                .writedata
			avs_cntl_byteenable  => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,              --                .byteenable
			avs_cntl_address     => "0"                                                                        --     (terminated)
		);

	ext_flash : component MebX_Qsys_Project_ext_flash
		generic map (
			TCM_ADDRESS_W                  => 26,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 100,
			TCM_WRITE_WAIT                 => 100,
			TCM_SETUP_WAIT                 => 25,
			TCM_DATA_HOLD                  => 20,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => m0_ddr3_memory_afi_half_clk_clk,               --   clk.clk
			reset_reset          => rst_controller_003_reset_out_reset,            -- reset.reset
			uas_address          => mm_interconnect_1_ext_flash_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_1_ext_flash_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_1_ext_flash_uas_read,          --      .read
			uas_write            => mm_interconnect_1_ext_flash_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_1_ext_flash_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_1_ext_flash_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_1_ext_flash_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_1_ext_flash_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_1_ext_flash_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_1_ext_flash_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_1_ext_flash_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ext_flash_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_n_out       => ext_flash_tcm_read_n_out,                      --      .read_n_out
			tcm_chipselect_n_out => ext_flash_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ext_flash_tcm_request,                         --      .request
			tcm_grant            => ext_flash_tcm_grant,                           --      .grant
			tcm_address_out      => ext_flash_tcm_address_out,                     --      .address_out
			tcm_data_out         => ext_flash_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ext_flash_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ext_flash_tcm_data_in                          --      .data_in
		);

	jtag_uart : component MebX_Qsys_Project_jtag_uart
		port map (
			clk            => m0_ddr3_memory_afi_half_clk_clk,                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	m0_ddr3_i2c_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m0_ddr3_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m0_ddr3_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m0_ddr3_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m0_ddr3_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m0_ddr3_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => m0_ddr3_i2c_scl_export                                -- external_connection.export
		);

	m0_ddr3_i2c_sda : component MebX_Qsys_Project_m0_ddr3_i2c_sda
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m0_ddr3_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m0_ddr3_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m0_ddr3_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m0_ddr3_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m0_ddr3_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => m0_ddr3_i2c_sda_export                                -- external_connection.export
		);

	m0_ddr3_memory : component MebX_Qsys_Project_m0_ddr3_memory
		port map (
			pll_ref_clk               => clk50_clk,                                               --      pll_ref_clk.clk
			global_reset_n            => rst_reset_n,                                             --     global_reset.reset_n
			soft_reset_n              => rst_reset_n,                                             --       soft_reset.reset_n
			afi_clk                   => m0_ddr3_memory_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk              => m0_ddr3_memory_afi_half_clk_clk,                         --     afi_half_clk.clk
			afi_reset_n               => open,                                                    --        afi_reset.reset_n
			afi_reset_export_n        => open,                                                    -- afi_reset_export.reset_n
			mem_a                     => m0_ddr3_memory_mem_a,                                    --           memory.mem_a
			mem_ba                    => m0_ddr3_memory_mem_ba,                                   --                 .mem_ba
			mem_ck                    => m0_ddr3_memory_mem_ck,                                   --                 .mem_ck
			mem_ck_n                  => m0_ddr3_memory_mem_ck_n,                                 --                 .mem_ck_n
			mem_cke                   => m0_ddr3_memory_mem_cke,                                  --                 .mem_cke
			mem_cs_n                  => m0_ddr3_memory_mem_cs_n,                                 --                 .mem_cs_n
			mem_dm                    => m0_ddr3_memory_mem_dm,                                   --                 .mem_dm
			mem_ras_n                 => m0_ddr3_memory_mem_ras_n,                                --                 .mem_ras_n
			mem_cas_n                 => m0_ddr3_memory_mem_cas_n,                                --                 .mem_cas_n
			mem_we_n                  => m0_ddr3_memory_mem_we_n,                                 --                 .mem_we_n
			mem_reset_n               => m0_ddr3_memory_mem_reset_n,                              --                 .mem_reset_n
			mem_dq                    => m0_ddr3_memory_mem_dq,                                   --                 .mem_dq
			mem_dqs                   => m0_ddr3_memory_mem_dqs,                                  --                 .mem_dqs
			mem_dqs_n                 => m0_ddr3_memory_mem_dqs_n,                                --                 .mem_dqs_n
			mem_odt                   => m0_ddr3_memory_mem_odt,                                  --                 .mem_odt
			avl_ready                 => m0_ddr3_memory_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin            => mm_interconnect_0_m0_ddr3_memory_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr                  => mm_interconnect_0_m0_ddr3_memory_avl_address,            --                 .address
			avl_rdata_valid           => mm_interconnect_0_m0_ddr3_memory_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata                 => mm_interconnect_0_m0_ddr3_memory_avl_readdata,           --                 .readdata
			avl_wdata                 => mm_interconnect_0_m0_ddr3_memory_avl_writedata,          --                 .writedata
			avl_be                    => mm_interconnect_0_m0_ddr3_memory_avl_byteenable,         --                 .byteenable
			avl_read_req              => mm_interconnect_0_m0_ddr3_memory_avl_read,               --                 .read
			avl_write_req             => mm_interconnect_0_m0_ddr3_memory_avl_write,              --                 .write
			avl_size                  => mm_interconnect_0_m0_ddr3_memory_avl_burstcount,         --                 .burstcount
			local_init_done           => m0_ddr3_memory_status_local_init_done,                   --           status.local_init_done
			local_cal_success         => m0_ddr3_memory_status_local_cal_success,                 --                 .local_cal_success
			local_cal_fail            => m0_ddr3_memory_status_local_cal_fail,                    --                 .local_cal_fail
			oct_rdn                   => m0_ddr3_oct_rdn,                                         --              oct.rdn
			oct_rup                   => m0_ddr3_oct_rup,                                         --                 .rup
			pll_mem_clk               => m0_ddr3_memory_pll_sharing_pll_mem_clk,                  --      pll_sharing.pll_mem_clk
			pll_write_clk             => m0_ddr3_memory_pll_sharing_pll_write_clk,                --                 .pll_write_clk
			pll_locked                => m0_ddr3_memory_pll_sharing_pll_locked,                   --                 .pll_locked
			pll_write_clk_pre_phy_clk => m0_ddr3_memory_pll_sharing_pll_write_clk_pre_phy_clk,    --                 .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          => m0_ddr3_memory_pll_sharing_pll_addr_cmd_clk,             --                 .pll_addr_cmd_clk
			pll_avl_clk               => m0_ddr3_memory_pll_sharing_pll_avl_clk,                  --                 .pll_avl_clk
			pll_config_clk            => m0_ddr3_memory_pll_sharing_pll_config_clk                --                 .pll_config_clk
		);

	nios2_gen2_0 : component MebX_Qsys_Project_nios2_gen2_0
		port map (
			clk                                 => m0_ddr3_memory_afi_half_clk_clk,                            --                       clk.clk
			reset_n                             => rst_controller_004_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_004_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_burstcount                        => nios2_gen2_0_instruction_master_burstcount,                 --                          .burstcount
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory : component MebX_Qsys_Project_onchip_memory
		port map (
			clk        => m0_ddr3_memory_afi_half_clk_clk,               --   clk1.clk
			address    => mm_interconnect_1_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_1_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_1_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	rst_controller : component rst_controller_top
		port map (
			clock_sink_clk                          => clk50_clk,                                                                --                  clock_sink.clk
			reset_sink_reset                        => rst_controller_002_reset_out_reset,                                       --                  reset_sink.reset
			reset_source_rs232_reset                => open,                                                                     --          reset_source_rs232.reset
			avalon_slave_rst_controller_address     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,     -- avalon_rst_controller_slave.address
			avalon_slave_rst_controller_write       => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,       --                            .write
			avalon_slave_rst_controller_read        => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,        --                            .read
			avalon_slave_rst_controller_writedata   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,   --                            .writedata
			avalon_slave_rst_controller_readdata    => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,    --                            .readdata
			avalon_slave_rst_controller_waitrequest => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest, --                            .waitrequest
			simucam_reset_signal                    => rst_controller_conduit_simucam_reset_t_simucam_reset_signal,              --       conduit_simucam_reset.t_simucam_reset_signal
			reset_input_signal                      => rst_controller_conduit_reset_input_t_reset_input_signal                   --         conduit_reset_input.t_reset_input_signal
		);

	sd_card_wp_n : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_sd_card_wp_n_s1_address,    --                  s1.address
			readdata => mm_interconnect_2_sd_card_wp_n_s1_readdata,   --                    .readdata
			in_port  => sd_card_wp_n_io_export                        -- external_connection.export
		);

	slide_sw : component MebX_Qsys_Project_button
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_002_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_slide_sw_s1_address,        --                  s1.address
			readdata => mm_interconnect_2_slide_sw_s1_readdata,       --                    .readdata
			in_port  => slide_sw_export                               -- external_connection.export
		);

	sysid_qsys : component MebX_Qsys_Project_sysid_qsys
		port map (
			clock    => m0_ddr3_memory_afi_half_clk_clk,                       --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	temp_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_scl_s1_readdata,        --                    .readdata
			out_port   => temp_scl_export                                -- external_connection.export
		);

	temp_sda : component MebX_Qsys_Project_m0_ddr3_i2c_sda
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_sda_s1_readdata,        --                    .readdata
			bidir_port => temp_sda_export                                -- external_connection.export
		);

	timer_1ms : component MebX_Qsys_Project_timer_1ms
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_002_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1ms_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1ms_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1ms_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1ms_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1ms_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_receiver_irq(0),               --           irq.irq
			timeout_pulse => timer_1ms_external_port_export                  -- external_port.export
		);

	timer_1us : component MebX_Qsys_Project_timer_1us
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_002_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1us_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1us_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1us_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1us_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1us_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_001_receiver_irq(0),           --           irq.irq
			timeout_pulse => timer_1us_external_port_export                  -- external_port.export
		);

	tristate_conduit_bridge_0 : component MebX_Qsys_Project_tristate_conduit_bridge_0
		port map (
			clk                         => m0_ddr3_memory_afi_half_clk_clk,       --   clk.clk
			reset                       => rst_controller_003_reset_out_reset,    -- reset.reset
			request                     => ext_flash_tcm_request,                 --   tcs.request
			grant                       => ext_flash_tcm_grant,                   --      .grant
			tcs_tcm_address_out         => ext_flash_tcm_address_out,             --      .address_out
			tcs_tcm_read_n_out(0)       => ext_flash_tcm_read_n_out,              --      .read_n_out
			tcs_tcm_write_n_out(0)      => ext_flash_tcm_write_n_out,             --      .write_n_out
			tcs_tcm_data_out            => ext_flash_tcm_data_out,                --      .data_out
			tcs_tcm_data_outen          => ext_flash_tcm_data_outen,              --      .data_outen
			tcs_tcm_data_in             => ext_flash_tcm_data_in,                 --      .data_in
			tcs_tcm_chipselect_n_out(0) => ext_flash_tcm_chipselect_n_out,        --      .chipselect_n_out
			tcm_address_out             => tristate_conduit_tcm_address_out,      --   out.tcm_address_out
			tcm_read_n_out              => tristate_conduit_tcm_read_n_out,       --      .tcm_read_n_out
			tcm_write_n_out             => tristate_conduit_tcm_write_n_out,      --      .tcm_write_n_out
			tcm_data_out                => tristate_conduit_tcm_data_out,         --      .tcm_data_out
			tcm_chipselect_n_out        => tristate_conduit_tcm_chipselect_n_out  --      .tcm_chipselect_n_out
		);

	mm_interconnect_0 : component MebX_Qsys_Project_mm_interconnect_0
		port map (
			clk_100_clk_clk                                                 => m0_ddr3_memory_afi_half_clk_clk,                          --                                               clk_100_clk.clk
			m0_ddr3_memory_afi_clk_clk                                      => m0_ddr3_memory_afi_clk_clk,                               --                                    m0_ddr3_memory_afi_clk.clk
			m0_ddr3_memory_avl_translator_reset_reset_bridge_in_reset_reset => rst_controller_005_reset_out_reset,                       -- m0_ddr3_memory_avl_translator_reset_reset_bridge_in_reset.reset
			m0_ddr3_memory_soft_reset_reset_bridge_in_reset_reset           => rst_controller_005_reset_out_reset,                       --           m0_ddr3_memory_soft_reset_reset_bridge_in_reset.reset
			Memory_Filler_reset_sink_reset_bridge_in_reset_reset            => rst_controller_001_reset_out_reset,                       --            Memory_Filler_reset_sink_reset_bridge_in_reset.reset
			ddr2_address_span_extender_expanded_master_address              => ddr2_address_span_extender_expanded_master_address,       --                ddr2_address_span_extender_expanded_master.address
			ddr2_address_span_extender_expanded_master_waitrequest          => ddr2_address_span_extender_expanded_master_waitrequest,   --                                                          .waitrequest
			ddr2_address_span_extender_expanded_master_burstcount           => ddr2_address_span_extender_expanded_master_burstcount,    --                                                          .burstcount
			ddr2_address_span_extender_expanded_master_byteenable           => ddr2_address_span_extender_expanded_master_byteenable,    --                                                          .byteenable
			ddr2_address_span_extender_expanded_master_read                 => ddr2_address_span_extender_expanded_master_read,          --                                                          .read
			ddr2_address_span_extender_expanded_master_readdata             => ddr2_address_span_extender_expanded_master_readdata,      --                                                          .readdata
			ddr2_address_span_extender_expanded_master_readdatavalid        => ddr2_address_span_extender_expanded_master_readdatavalid, --                                                          .readdatavalid
			ddr2_address_span_extender_expanded_master_write                => ddr2_address_span_extender_expanded_master_write,         --                                                          .write
			ddr2_address_span_extender_expanded_master_writedata            => ddr2_address_span_extender_expanded_master_writedata,     --                                                          .writedata
			Memory_Filler_avalon_master_data_address                        => memory_filler_avalon_master_data_address,                 --                          Memory_Filler_avalon_master_data.address
			Memory_Filler_avalon_master_data_waitrequest                    => memory_filler_avalon_master_data_waitrequest,             --                                                          .waitrequest
			Memory_Filler_avalon_master_data_write                          => memory_filler_avalon_master_data_write,                   --                                                          .write
			Memory_Filler_avalon_master_data_writedata                      => memory_filler_avalon_master_data_writedata,               --                                                          .writedata
			m0_ddr3_memory_avl_address                                      => mm_interconnect_0_m0_ddr3_memory_avl_address,             --                                        m0_ddr3_memory_avl.address
			m0_ddr3_memory_avl_write                                        => mm_interconnect_0_m0_ddr3_memory_avl_write,               --                                                          .write
			m0_ddr3_memory_avl_read                                         => mm_interconnect_0_m0_ddr3_memory_avl_read,                --                                                          .read
			m0_ddr3_memory_avl_readdata                                     => mm_interconnect_0_m0_ddr3_memory_avl_readdata,            --                                                          .readdata
			m0_ddr3_memory_avl_writedata                                    => mm_interconnect_0_m0_ddr3_memory_avl_writedata,           --                                                          .writedata
			m0_ddr3_memory_avl_beginbursttransfer                           => mm_interconnect_0_m0_ddr3_memory_avl_beginbursttransfer,  --                                                          .beginbursttransfer
			m0_ddr3_memory_avl_burstcount                                   => mm_interconnect_0_m0_ddr3_memory_avl_burstcount,          --                                                          .burstcount
			m0_ddr3_memory_avl_byteenable                                   => mm_interconnect_0_m0_ddr3_memory_avl_byteenable,          --                                                          .byteenable
			m0_ddr3_memory_avl_readdatavalid                                => mm_interconnect_0_m0_ddr3_memory_avl_readdatavalid,       --                                                          .readdatavalid
			m0_ddr3_memory_avl_waitrequest                                  => mm_interconnect_0_m0_ddr3_memory_avl_inv                  --                                                          .waitrequest
		);

	mm_interconnect_1 : component MebX_Qsys_Project_mm_interconnect_1
		port map (
			clk_100_clk_clk                                         => m0_ddr3_memory_afi_half_clk_clk,                                           --                               clk_100_clk.clk
			ext_flash_reset_reset_bridge_in_reset_reset             => rst_controller_003_reset_out_reset,                                        --     ext_flash_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset             => rst_controller_001_reset_out_reset,                                        --     jtag_uart_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset          => rst_controller_004_reset_out_reset,                                        --  nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                        => nios2_gen2_0_data_master_address,                                          --                  nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                    => nios2_gen2_0_data_master_waitrequest,                                      --                                          .waitrequest
			nios2_gen2_0_data_master_byteenable                     => nios2_gen2_0_data_master_byteenable,                                       --                                          .byteenable
			nios2_gen2_0_data_master_read                           => nios2_gen2_0_data_master_read,                                             --                                          .read
			nios2_gen2_0_data_master_readdata                       => nios2_gen2_0_data_master_readdata,                                         --                                          .readdata
			nios2_gen2_0_data_master_write                          => nios2_gen2_0_data_master_write,                                            --                                          .write
			nios2_gen2_0_data_master_writedata                      => nios2_gen2_0_data_master_writedata,                                        --                                          .writedata
			nios2_gen2_0_data_master_debugaccess                    => nios2_gen2_0_data_master_debugaccess,                                      --                                          .debugaccess
			nios2_gen2_0_instruction_master_address                 => nios2_gen2_0_instruction_master_address,                                   --           nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest             => nios2_gen2_0_instruction_master_waitrequest,                               --                                          .waitrequest
			nios2_gen2_0_instruction_master_burstcount              => nios2_gen2_0_instruction_master_burstcount,                                --                                          .burstcount
			nios2_gen2_0_instruction_master_read                    => nios2_gen2_0_instruction_master_read,                                      --                                          .read
			nios2_gen2_0_instruction_master_readdata                => nios2_gen2_0_instruction_master_readdata,                                  --                                          .readdata
			nios2_gen2_0_instruction_master_readdatavalid           => nios2_gen2_0_instruction_master_readdatavalid,                             --                                          .readdatavalid
			clock_bridge_afi_50_s0_address                          => mm_interconnect_1_clock_bridge_afi_50_s0_address,                          --                    clock_bridge_afi_50_s0.address
			clock_bridge_afi_50_s0_write                            => mm_interconnect_1_clock_bridge_afi_50_s0_write,                            --                                          .write
			clock_bridge_afi_50_s0_read                             => mm_interconnect_1_clock_bridge_afi_50_s0_read,                             --                                          .read
			clock_bridge_afi_50_s0_readdata                         => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,                         --                                          .readdata
			clock_bridge_afi_50_s0_writedata                        => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,                        --                                          .writedata
			clock_bridge_afi_50_s0_burstcount                       => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,                       --                                          .burstcount
			clock_bridge_afi_50_s0_byteenable                       => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,                       --                                          .byteenable
			clock_bridge_afi_50_s0_readdatavalid                    => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid,                    --                                          .readdatavalid
			clock_bridge_afi_50_s0_waitrequest                      => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,                      --                                          .waitrequest
			clock_bridge_afi_50_s0_debugaccess                      => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,                      --                                          .debugaccess
			ddr2_address_span_extender_cntl_write                   => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                   --           ddr2_address_span_extender_cntl.write
			ddr2_address_span_extender_cntl_read                    => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                    --                                          .read
			ddr2_address_span_extender_cntl_readdata                => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                --                                          .readdata
			ddr2_address_span_extender_cntl_writedata               => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,               --                                          .writedata
			ddr2_address_span_extender_cntl_byteenable              => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,              --                                          .byteenable
			ddr2_address_span_extender_windowed_slave_address       => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,       -- ddr2_address_span_extender_windowed_slave.address
			ddr2_address_span_extender_windowed_slave_write         => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,         --                                          .write
			ddr2_address_span_extender_windowed_slave_read          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,          --                                          .read
			ddr2_address_span_extender_windowed_slave_readdata      => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,      --                                          .readdata
			ddr2_address_span_extender_windowed_slave_writedata     => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,     --                                          .writedata
			ddr2_address_span_extender_windowed_slave_burstcount    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,    --                                          .burstcount
			ddr2_address_span_extender_windowed_slave_byteenable    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,    --                                          .byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid, --                                          .readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest   => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,   --                                          .waitrequest
			ext_flash_uas_address                                   => mm_interconnect_1_ext_flash_uas_address,                                   --                             ext_flash_uas.address
			ext_flash_uas_write                                     => mm_interconnect_1_ext_flash_uas_write,                                     --                                          .write
			ext_flash_uas_read                                      => mm_interconnect_1_ext_flash_uas_read,                                      --                                          .read
			ext_flash_uas_readdata                                  => mm_interconnect_1_ext_flash_uas_readdata,                                  --                                          .readdata
			ext_flash_uas_writedata                                 => mm_interconnect_1_ext_flash_uas_writedata,                                 --                                          .writedata
			ext_flash_uas_burstcount                                => mm_interconnect_1_ext_flash_uas_burstcount,                                --                                          .burstcount
			ext_flash_uas_byteenable                                => mm_interconnect_1_ext_flash_uas_byteenable,                                --                                          .byteenable
			ext_flash_uas_readdatavalid                             => mm_interconnect_1_ext_flash_uas_readdatavalid,                             --                                          .readdatavalid
			ext_flash_uas_waitrequest                               => mm_interconnect_1_ext_flash_uas_waitrequest,                               --                                          .waitrequest
			ext_flash_uas_lock                                      => mm_interconnect_1_ext_flash_uas_lock,                                      --                                          .lock
			ext_flash_uas_debugaccess                               => mm_interconnect_1_ext_flash_uas_debugaccess,                               --                                          .debugaccess
			jtag_uart_avalon_jtag_slave_address                     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,                     --               jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                       => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,                       --                                          .write
			jtag_uart_avalon_jtag_slave_read                        => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,                        --                                          .read
			jtag_uart_avalon_jtag_slave_readdata                    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,                    --                                          .readdata
			jtag_uart_avalon_jtag_slave_writedata                   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,                   --                                          .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                 => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,                 --                                          .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,                  --                                          .chipselect
			Memory_Filler_avalon_slave_config_address               => mm_interconnect_1_memory_filler_avalon_slave_config_address,               --         Memory_Filler_avalon_slave_config.address
			Memory_Filler_avalon_slave_config_write                 => mm_interconnect_1_memory_filler_avalon_slave_config_write,                 --                                          .write
			Memory_Filler_avalon_slave_config_read                  => mm_interconnect_1_memory_filler_avalon_slave_config_read,                  --                                          .read
			Memory_Filler_avalon_slave_config_readdata              => mm_interconnect_1_memory_filler_avalon_slave_config_readdata,              --                                          .readdata
			Memory_Filler_avalon_slave_config_writedata             => mm_interconnect_1_memory_filler_avalon_slave_config_writedata,             --                                          .writedata
			Memory_Filler_avalon_slave_config_byteenable            => mm_interconnect_1_memory_filler_avalon_slave_config_byteenable,            --                                          .byteenable
			Memory_Filler_avalon_slave_config_waitrequest           => mm_interconnect_1_memory_filler_avalon_slave_config_waitrequest,           --                                          .waitrequest
			nios2_gen2_0_debug_mem_slave_address                    => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,                    --              nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                      => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,                      --                                          .write
			nios2_gen2_0_debug_mem_slave_read                       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,                       --                                          .read
			nios2_gen2_0_debug_mem_slave_readdata                   => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,                   --                                          .readdata
			nios2_gen2_0_debug_mem_slave_writedata                  => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,                  --                                          .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                 => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,                 --                                          .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest,                --                                          .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess,                --                                          .debugaccess
			onchip_memory_s1_address                                => mm_interconnect_1_onchip_memory_s1_address,                                --                          onchip_memory_s1.address
			onchip_memory_s1_write                                  => mm_interconnect_1_onchip_memory_s1_write,                                  --                                          .write
			onchip_memory_s1_readdata                               => mm_interconnect_1_onchip_memory_s1_readdata,                               --                                          .readdata
			onchip_memory_s1_writedata                              => mm_interconnect_1_onchip_memory_s1_writedata,                              --                                          .writedata
			onchip_memory_s1_byteenable                             => mm_interconnect_1_onchip_memory_s1_byteenable,                             --                                          .byteenable
			onchip_memory_s1_chipselect                             => mm_interconnect_1_onchip_memory_s1_chipselect,                             --                                          .chipselect
			onchip_memory_s1_clken                                  => mm_interconnect_1_onchip_memory_s1_clken,                                  --                                          .clken
			sysid_qsys_control_slave_address                        => mm_interconnect_1_sysid_qsys_control_slave_address,                        --                  sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                       => mm_interconnect_1_sysid_qsys_control_slave_readdata                        --                                          .readdata
		);

	mm_interconnect_2 : component MebX_Qsys_Project_mm_interconnect_2
		port map (
			clk_50_clk_clk                                           => clk50_clk,                                                                --                                         clk_50_clk.clk
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                       -- clock_bridge_afi_50_m0_reset_reset_bridge_in_reset.reset
			clock_bridge_afi_50_m0_address                           => clock_bridge_afi_50_m0_address,                                           --                             clock_bridge_afi_50_m0.address
			clock_bridge_afi_50_m0_waitrequest                       => clock_bridge_afi_50_m0_waitrequest,                                       --                                                   .waitrequest
			clock_bridge_afi_50_m0_burstcount                        => clock_bridge_afi_50_m0_burstcount,                                        --                                                   .burstcount
			clock_bridge_afi_50_m0_byteenable                        => clock_bridge_afi_50_m0_byteenable,                                        --                                                   .byteenable
			clock_bridge_afi_50_m0_read                              => clock_bridge_afi_50_m0_read,                                              --                                                   .read
			clock_bridge_afi_50_m0_readdata                          => clock_bridge_afi_50_m0_readdata,                                          --                                                   .readdata
			clock_bridge_afi_50_m0_readdatavalid                     => clock_bridge_afi_50_m0_readdatavalid,                                     --                                                   .readdatavalid
			clock_bridge_afi_50_m0_write                             => clock_bridge_afi_50_m0_write,                                             --                                                   .write
			clock_bridge_afi_50_m0_writedata                         => clock_bridge_afi_50_m0_writedata,                                         --                                                   .writedata
			clock_bridge_afi_50_m0_debugaccess                       => clock_bridge_afi_50_m0_debugaccess,                                       --                                                   .debugaccess
			board_led_s1_address                                     => mm_interconnect_2_board_led_s1_address,                                   --                                       board_led_s1.address
			board_led_s1_write                                       => mm_interconnect_2_board_led_s1_write,                                     --                                                   .write
			board_led_s1_readdata                                    => mm_interconnect_2_board_led_s1_readdata,                                  --                                                   .readdata
			board_led_s1_writedata                                   => mm_interconnect_2_board_led_s1_writedata,                                 --                                                   .writedata
			board_led_s1_chipselect                                  => mm_interconnect_2_board_led_s1_chipselect,                                --                                                   .chipselect
			button_s1_address                                        => mm_interconnect_2_button_s1_address,                                      --                                          button_s1.address
			button_s1_readdata                                       => mm_interconnect_2_button_s1_readdata,                                     --                                                   .readdata
			csense_adc_fo_s1_address                                 => mm_interconnect_2_csense_adc_fo_s1_address,                               --                                   csense_adc_fo_s1.address
			csense_adc_fo_s1_write                                   => mm_interconnect_2_csense_adc_fo_s1_write,                                 --                                                   .write
			csense_adc_fo_s1_readdata                                => mm_interconnect_2_csense_adc_fo_s1_readdata,                              --                                                   .readdata
			csense_adc_fo_s1_writedata                               => mm_interconnect_2_csense_adc_fo_s1_writedata,                             --                                                   .writedata
			csense_adc_fo_s1_chipselect                              => mm_interconnect_2_csense_adc_fo_s1_chipselect,                            --                                                   .chipselect
			csense_cs_n_s1_address                                   => mm_interconnect_2_csense_cs_n_s1_address,                                 --                                     csense_cs_n_s1.address
			csense_cs_n_s1_write                                     => mm_interconnect_2_csense_cs_n_s1_write,                                   --                                                   .write
			csense_cs_n_s1_readdata                                  => mm_interconnect_2_csense_cs_n_s1_readdata,                                --                                                   .readdata
			csense_cs_n_s1_writedata                                 => mm_interconnect_2_csense_cs_n_s1_writedata,                               --                                                   .writedata
			csense_cs_n_s1_chipselect                                => mm_interconnect_2_csense_cs_n_s1_chipselect,                              --                                                   .chipselect
			csense_sck_s1_address                                    => mm_interconnect_2_csense_sck_s1_address,                                  --                                      csense_sck_s1.address
			csense_sck_s1_write                                      => mm_interconnect_2_csense_sck_s1_write,                                    --                                                   .write
			csense_sck_s1_readdata                                   => mm_interconnect_2_csense_sck_s1_readdata,                                 --                                                   .readdata
			csense_sck_s1_writedata                                  => mm_interconnect_2_csense_sck_s1_writedata,                                --                                                   .writedata
			csense_sck_s1_chipselect                                 => mm_interconnect_2_csense_sck_s1_chipselect,                               --                                                   .chipselect
			csense_sdi_s1_address                                    => mm_interconnect_2_csense_sdi_s1_address,                                  --                                      csense_sdi_s1.address
			csense_sdi_s1_write                                      => mm_interconnect_2_csense_sdi_s1_write,                                    --                                                   .write
			csense_sdi_s1_readdata                                   => mm_interconnect_2_csense_sdi_s1_readdata,                                 --                                                   .readdata
			csense_sdi_s1_writedata                                  => mm_interconnect_2_csense_sdi_s1_writedata,                                --                                                   .writedata
			csense_sdi_s1_chipselect                                 => mm_interconnect_2_csense_sdi_s1_chipselect,                               --                                                   .chipselect
			csense_sdo_s1_address                                    => mm_interconnect_2_csense_sdo_s1_address,                                  --                                      csense_sdo_s1.address
			csense_sdo_s1_readdata                                   => mm_interconnect_2_csense_sdo_s1_readdata,                                 --                                                   .readdata
			m0_ddr3_i2c_scl_s1_address                               => mm_interconnect_2_m0_ddr3_i2c_scl_s1_address,                             --                                 m0_ddr3_i2c_scl_s1.address
			m0_ddr3_i2c_scl_s1_write                                 => mm_interconnect_2_m0_ddr3_i2c_scl_s1_write,                               --                                                   .write
			m0_ddr3_i2c_scl_s1_readdata                              => mm_interconnect_2_m0_ddr3_i2c_scl_s1_readdata,                            --                                                   .readdata
			m0_ddr3_i2c_scl_s1_writedata                             => mm_interconnect_2_m0_ddr3_i2c_scl_s1_writedata,                           --                                                   .writedata
			m0_ddr3_i2c_scl_s1_chipselect                            => mm_interconnect_2_m0_ddr3_i2c_scl_s1_chipselect,                          --                                                   .chipselect
			m0_ddr3_i2c_sda_s1_address                               => mm_interconnect_2_m0_ddr3_i2c_sda_s1_address,                             --                                 m0_ddr3_i2c_sda_s1.address
			m0_ddr3_i2c_sda_s1_write                                 => mm_interconnect_2_m0_ddr3_i2c_sda_s1_write,                               --                                                   .write
			m0_ddr3_i2c_sda_s1_readdata                              => mm_interconnect_2_m0_ddr3_i2c_sda_s1_readdata,                            --                                                   .readdata
			m0_ddr3_i2c_sda_s1_writedata                             => mm_interconnect_2_m0_ddr3_i2c_sda_s1_writedata,                           --                                                   .writedata
			m0_ddr3_i2c_sda_s1_chipselect                            => mm_interconnect_2_m0_ddr3_i2c_sda_s1_chipselect,                          --                                                   .chipselect
			rst_controller_avalon_rst_controller_slave_address       => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,     --         rst_controller_avalon_rst_controller_slave.address
			rst_controller_avalon_rst_controller_slave_write         => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,       --                                                   .write
			rst_controller_avalon_rst_controller_slave_read          => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,        --                                                   .read
			rst_controller_avalon_rst_controller_slave_readdata      => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,    --                                                   .readdata
			rst_controller_avalon_rst_controller_slave_writedata     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,   --                                                   .writedata
			rst_controller_avalon_rst_controller_slave_waitrequest   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest, --                                                   .waitrequest
			sd_card_wp_n_s1_address                                  => mm_interconnect_2_sd_card_wp_n_s1_address,                                --                                    sd_card_wp_n_s1.address
			sd_card_wp_n_s1_readdata                                 => mm_interconnect_2_sd_card_wp_n_s1_readdata,                               --                                                   .readdata
			slide_sw_s1_address                                      => mm_interconnect_2_slide_sw_s1_address,                                    --                                        slide_sw_s1.address
			slide_sw_s1_readdata                                     => mm_interconnect_2_slide_sw_s1_readdata,                                   --                                                   .readdata
			temp_scl_s1_address                                      => mm_interconnect_2_temp_scl_s1_address,                                    --                                        temp_scl_s1.address
			temp_scl_s1_write                                        => mm_interconnect_2_temp_scl_s1_write,                                      --                                                   .write
			temp_scl_s1_readdata                                     => mm_interconnect_2_temp_scl_s1_readdata,                                   --                                                   .readdata
			temp_scl_s1_writedata                                    => mm_interconnect_2_temp_scl_s1_writedata,                                  --                                                   .writedata
			temp_scl_s1_chipselect                                   => mm_interconnect_2_temp_scl_s1_chipselect,                                 --                                                   .chipselect
			temp_sda_s1_address                                      => mm_interconnect_2_temp_sda_s1_address,                                    --                                        temp_sda_s1.address
			temp_sda_s1_write                                        => mm_interconnect_2_temp_sda_s1_write,                                      --                                                   .write
			temp_sda_s1_readdata                                     => mm_interconnect_2_temp_sda_s1_readdata,                                   --                                                   .readdata
			temp_sda_s1_writedata                                    => mm_interconnect_2_temp_sda_s1_writedata,                                  --                                                   .writedata
			temp_sda_s1_chipselect                                   => mm_interconnect_2_temp_sda_s1_chipselect,                                 --                                                   .chipselect
			timer_1ms_s1_address                                     => mm_interconnect_2_timer_1ms_s1_address,                                   --                                       timer_1ms_s1.address
			timer_1ms_s1_write                                       => mm_interconnect_2_timer_1ms_s1_write,                                     --                                                   .write
			timer_1ms_s1_readdata                                    => mm_interconnect_2_timer_1ms_s1_readdata,                                  --                                                   .readdata
			timer_1ms_s1_writedata                                   => mm_interconnect_2_timer_1ms_s1_writedata,                                 --                                                   .writedata
			timer_1ms_s1_chipselect                                  => mm_interconnect_2_timer_1ms_s1_chipselect,                                --                                                   .chipselect
			timer_1us_s1_address                                     => mm_interconnect_2_timer_1us_s1_address,                                   --                                       timer_1us_s1.address
			timer_1us_s1_write                                       => mm_interconnect_2_timer_1us_s1_write,                                     --                                                   .write
			timer_1us_s1_readdata                                    => mm_interconnect_2_timer_1us_s1_readdata,                                  --                                                   .readdata
			timer_1us_s1_writedata                                   => mm_interconnect_2_timer_1us_s1_writedata,                                 --                                                   .writedata
			timer_1us_s1_chipselect                                  => mm_interconnect_2_timer_1us_s1_chipselect                                 --                                                   .chipselect
		);

	irq_mapper : component MebX_Qsys_Project_irq_mapper
		port map (
			clk           => m0_ddr3_memory_afi_half_clk_clk,    --       clk.clk
			reset         => rst_controller_004_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m0_ddr3_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_002_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_004_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m0_ddr3_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_002_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_004_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	rst_controller_001 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m0_ddr3_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component mebx_qsys_project_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => clk50_clk,                          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component mebx_qsys_project_rst_controller_003
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => rst_reset_n_ports_inv,              -- reset_in1.reset
			clk            => m0_ddr3_memory_afi_half_clk_clk,    --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m0_ddr3_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_004_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_005 : component mebx_qsys_project_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m0_ddr3_memory_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_reset_n_ports_inv <= not rst_reset_n;

	mm_interconnect_0_m0_ddr3_memory_avl_inv <= not m0_ddr3_memory_avl_waitrequest;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_2_timer_1ms_s1_write_ports_inv <= not mm_interconnect_2_timer_1ms_s1_write;

	mm_interconnect_2_timer_1us_s1_write_ports_inv <= not mm_interconnect_2_timer_1us_s1_write;

	mm_interconnect_2_temp_scl_s1_write_ports_inv <= not mm_interconnect_2_temp_scl_s1_write;

	mm_interconnect_2_temp_sda_s1_write_ports_inv <= not mm_interconnect_2_temp_sda_s1_write;

	mm_interconnect_2_m0_ddr3_i2c_sda_s1_write_ports_inv <= not mm_interconnect_2_m0_ddr3_i2c_sda_s1_write;

	mm_interconnect_2_m0_ddr3_i2c_scl_s1_write_ports_inv <= not mm_interconnect_2_m0_ddr3_i2c_scl_s1_write;

	mm_interconnect_2_csense_sdi_s1_write_ports_inv <= not mm_interconnect_2_csense_sdi_s1_write;

	mm_interconnect_2_csense_sck_s1_write_ports_inv <= not mm_interconnect_2_csense_sck_s1_write;

	mm_interconnect_2_csense_cs_n_s1_write_ports_inv <= not mm_interconnect_2_csense_cs_n_s1_write;

	mm_interconnect_2_csense_adc_fo_s1_write_ports_inv <= not mm_interconnect_2_csense_adc_fo_s1_write;

	mm_interconnect_2_board_led_s1_write_ports_inv <= not mm_interconnect_2_board_led_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

end architecture rtl; -- of MebX_Qsys_Project
